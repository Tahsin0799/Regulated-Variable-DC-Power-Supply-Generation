* E:\OneDrive - BUET\Tahsin\CODING ZONE\PSPICE Simulation\ALL EXPERIMENTS\EEE 208\OP-AMP\Regulated Variable DC Power Supply Generation\Final_ckt.sch

* Schematics Version 9.2
* Tue Feb 22 16:11:07 2022


.PARAM         var1=1k 

** Analysis setup **
.tran 30u 0.28 0 30u
.STEP LIN PARAM var1 50 3k 100 
.OP 


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "Final_ckt.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
