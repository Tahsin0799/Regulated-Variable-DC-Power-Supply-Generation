* E:\OneDrive - BUET\Tahsin\CODING ZONE\PSPICE Simulation\ALL EXPERIMENTS\EEE 208\OP-AMP\Regulated Variable DC Power Supply Generation\Regulation_process.sch

* Schematics Version 9.2
* Sun Feb 20 17:55:19 2022



** Analysis setup **
.tran 30u 0.28 0 30u
.OP 


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "Regulation_process.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
